module XSTop_wrapper(
  input           sys_clk_i,    
  input           sys_rstn_i, 
  input           osc_clock,        //24MHz
  input           outer_clock,      //Max : 2.4GHz
  input           global_reset,     //24MHz
  input           rtc_clk,          //1MHz

  input  [3:0]    pll_bypass_sel,   //apb clk : 100MHz
  output          pll0_lock,
  output          pll0_clk_div_1024,
  output [11:0]   pll0_test_calout,

  input  [15:0]   soc_to_cpu,   // none
  output [15:0]   cpu_to_soc,   //none

  input  [63:0]   io_extIntrs,   // come from IPs, Max : 600MHz

  input  [15:0]   io_sram_config,  //apb clk : 100MHz

  input           io_systemjtag_jtag_TCK,         // come from gpio
  input           io_systemjtag_jtag_TMS,         // come from gpio
  input           io_systemjtag_jtag_TDI,         // come from gpio
  output          io_systemjtag_jtag_TDO_data,    // come from gpio
  output          io_systemjtag_jtag_TDO_driven,  // come from gpio
  input           io_systemjtag_reset,            // come from gpio

// peri bus   //400MHz
// dma bus    //800MHz
// mem bus    //800MHz

  (*mark_debug="true"*) output          dma_core_awready,
  (*mark_debug="true"*) input           dma_core_awvalid,
  (*mark_debug="true"*) input  [13:0]   dma_core_awid,
  (*mark_debug="true"*) input  [35:0]   dma_core_awaddr,
  (*mark_debug="true"*) input  [7:0]    dma_core_awlen,
  (*mark_debug="true"*) input  [2:0]    dma_core_awsize,
  (*mark_debug="true"*) input  [1:0]    dma_core_awburst,
  (*mark_debug="true"*) input           dma_core_awlock,
  (*mark_debug="true"*) input  [3:0]    dma_core_awcache,
  (*mark_debug="true"*) input  [2:0]    dma_core_awprot,
  (*mark_debug="true"*) input  [3:0]    dma_core_awqos,
  (*mark_debug="true"*) output          dma_core_wready,
  (*mark_debug="true"*) input           dma_core_wvalid,
  (*mark_debug="true"*) input  [255:0]  dma_core_wdata,
  (*mark_debug="true"*) input  [31:0]   dma_core_wstrb,
  (*mark_debug="true"*) input           dma_core_wlast,
  (*mark_debug="true"*) input           dma_core_bready,
  (*mark_debug="true"*) output          dma_core_bvalid,
  (*mark_debug="true"*) output [13:0]   dma_core_bid,
  (*mark_debug="true"*) output [1:0]    dma_core_bresp,
  (*mark_debug="true"*) output          dma_core_arready,
  (*mark_debug="true"*) input           dma_core_arvalid,
  (*mark_debug="true"*) input  [13:0]   dma_core_arid,
  (*mark_debug="true"*) input  [35:0]   dma_core_araddr,
  (*mark_debug="true"*) input  [7:0]    dma_core_arlen,
  (*mark_debug="true"*) input  [2:0]    dma_core_arsize,
  (*mark_debug="true"*) input  [1:0]    dma_core_arburst,
  (*mark_debug="true"*) input           dma_core_arlock,
  (*mark_debug="true"*) input  [3:0]    dma_core_arcache,
  (*mark_debug="true"*) input  [2:0]    dma_core_arprot,
  (*mark_debug="true"*) input  [3:0]    dma_core_arqos,
  (*mark_debug="true"*) input           dma_core_rready,
  (*mark_debug="true"*) output          dma_core_rvalid,
  (*mark_debug="true"*) output [13:0]   dma_core_rid,
  (*mark_debug="true"*) output [255:0]  dma_core_rdata,
  (*mark_debug="true"*) output [1:0]    dma_core_rresp,
  (*mark_debug="true"*) output          dma_core_rlast,
  
  (*mark_debug="true"*) input           peri_awready,
  (*mark_debug="true"*) output          peri_awvalid,
  (*mark_debug="true"*) output [1:0]    peri_awid,
  (*mark_debug="true"*) output [30:0]   peri_awaddr,
  (*mark_debug="true"*) output [7:0]    peri_awlen,
  (*mark_debug="true"*) output [2:0]    peri_awsize,
  (*mark_debug="true"*) output [1:0]    peri_awburst,
  (*mark_debug="true"*) output          peri_awlock,
  (*mark_debug="true"*) output [3:0]    peri_awcache,
  (*mark_debug="true"*) output [2:0]    peri_awprot,
  (*mark_debug="true"*) output [3:0]    peri_awqos,
  (*mark_debug="true"*) input           peri_wready,
  (*mark_debug="true"*) output          peri_wvalid,
  (*mark_debug="true"*) output [63:0]   peri_wdata,
  (*mark_debug="true"*) output [7:0]    peri_wstrb,
  (*mark_debug="true"*) output          peri_wlast,
  (*mark_debug="true"*) output          peri_bready,
  (*mark_debug="true"*) input           peri_bvalid,
  (*mark_debug="true"*) input  [1:0]    peri_bid,
  (*mark_debug="true"*) input  [1:0]    peri_bresp,
  (*mark_debug="true"*) input           peri_arready,
  (*mark_debug="true"*) output          peri_arvalid,
  (*mark_debug="true"*) output [1:0]    peri_arid,
  (*mark_debug="true"*) output [30:0]   peri_araddr,
  (*mark_debug="true"*) output [7:0]    peri_arlen,
  (*mark_debug="true"*) output [2:0]    peri_arsize,
  (*mark_debug="true"*) output [1:0]    peri_arburst,
  (*mark_debug="true"*) output          peri_arlock,
  (*mark_debug="true"*) output [3:0]    peri_arcache,
  (*mark_debug="true"*) output [2:0]    peri_arprot,
  (*mark_debug="true"*) output [3:0]    peri_arqos,
  (*mark_debug="true"*) output          peri_rready,
  (*mark_debug="true"*) input           peri_rvalid,
  (*mark_debug="true"*) input  [1:0]    peri_rid,
  (*mark_debug="true"*) input  [63:0]   peri_rdata,
  (*mark_debug="true"*) input  [1:0]    peri_rresp,
  (*mark_debug="true"*) input           peri_rlast,
  
  (*mark_debug="true"*) input           mem_core_awready,
  (*mark_debug="true"*) output          mem_core_awvalid,
  (*mark_debug="true"*) output [13:0]   mem_core_awid,
  (*mark_debug="true"*) output [35:0]   mem_core_awaddr,
  (*mark_debug="true"*) output [7:0]    mem_core_awlen,
  (*mark_debug="true"*) output [2:0]    mem_core_awsize,
  (*mark_debug="true"*) output [1:0]    mem_core_awburst,
  (*mark_debug="true"*) output          mem_core_awlock,
  (*mark_debug="true"*) output [3:0]    mem_core_awcache,
  (*mark_debug="true"*) output [2:0]    mem_core_awprot,
  (*mark_debug="true"*) output [3:0]    mem_core_awqos,
  (*mark_debug="true"*) input           mem_core_wready,
  (*mark_debug="true"*) output          mem_core_wvalid,
  (*mark_debug="true"*) output [255:0]  mem_core_wdata,
  (*mark_debug="true"*) output [31:0]   mem_core_wstrb,
  (*mark_debug="true"*) output          mem_core_wlast,
  (*mark_debug="true"*) output          mem_core_bready,
  (*mark_debug="true"*) input           mem_core_bvalid,
  (*mark_debug="true"*) input  [13:0]   mem_core_bid,
  (*mark_debug="true"*) input  [1:0]    mem_core_bresp,
  (*mark_debug="true"*) input           mem_core_arready,
  (*mark_debug="true"*) output          mem_core_arvalid,
  (*mark_debug="true"*) output [13:0]   mem_core_arid,
  (*mark_debug="true"*) output [35:0]   mem_core_araddr,
  (*mark_debug="true"*) output [7:0]    mem_core_arlen,
  (*mark_debug="true"*) output [2:0]    mem_core_arsize,
  (*mark_debug="true"*) output [1:0]    mem_core_arburst,
  (*mark_debug="true"*) output          mem_core_arlock,
  (*mark_debug="true"*) output [3:0]    mem_core_arcache,
  (*mark_debug="true"*) output [2:0]    mem_core_arprot,
  (*mark_debug="true"*) output [3:0]    mem_core_arqos,
  (*mark_debug="true"*) output          mem_core_rready,
  (*mark_debug="true"*) input           mem_core_rvalid,
  (*mark_debug="true"*) input  [13:0]   mem_core_rid,
  (*mark_debug="true"*) input  [255:0]  mem_core_rdata,
  (*mark_debug="true"*) input  [1:0]    mem_core_rresp,
  (*mark_debug="true"*) input           mem_core_rlast
);

  wire          cpu_clock       ;
  wire          cpu_global_reset;
  wire          global_reset_sync;

  wire [31:0]   pll0_config_0;
  wire [31:0]   pll0_config_1;
  wire [31:0]   pll0_config_2;
  wire [31:0]   pll0_config_3;
  wire [31:0]   pll0_config_4;
  wire [31:0]   pll0_config_5;
//  wire [31:0]   pll0_config_5 = 32'h3;

assign cpu_to_soc = 32'h0;


XSTop  u_XSTop(
.m_memory_aw_ready                (mem_core_awready )                        ,
  .m_memory_aw_valid                (mem_core_awvalid )                        ,
  .m_memory_aw_id                  (mem_core_awid    )                          ,
  .m_memory_aw_addr                (mem_core_awaddr  )                            ,
  .m_memory_aw_len                 (mem_core_awlen   )                           ,
  .m_memory_aw_size                (mem_core_awsize  )                            ,
  .m_memory_aw_burst                (mem_core_awburst )                             ,
  .m_memory_aw_lock                (mem_core_awlock  )                            ,
  .m_memory_aw_cache                (mem_core_awcache )                             ,
  .m_memory_aw_prot                (mem_core_awprot  )                            ,
  .m_memory_aw_qos                 (mem_core_awqos   )                           ,
  .m_memory_w_ready                (mem_core_wready  )                       ,
  .m_memory_w_valid                (mem_core_wvalid  )                       ,
  .m_memory_w_data                 (mem_core_wdata   )                           ,
  .m_memory_w_strb                 (mem_core_wstrb   )                           ,
  .m_memory_w_last                 (mem_core_wlast   )                           ,
  .m_memory_b_ready                (mem_core_bready  )                       ,
  .m_memory_b_valid                (mem_core_bvalid  )                       ,
  .m_memory_b_id                   (mem_core_bid     )                         ,
  .m_memory_b_resp                 (mem_core_bresp   )                           ,
  .m_memory_ar_ready               (mem_core_arready )                        ,
  .m_memory_ar_valid                (mem_core_arvalid )                        ,
  .m_memory_ar_id                  (mem_core_arid    )                          ,
  .m_memory_ar_addr                (mem_core_araddr  )                            ,
  .m_memory_ar_len                 (mem_core_arlen   )                           ,
  .m_memory_ar_size                (mem_core_arsize  )                            ,
  .m_memory_ar_burst                (mem_core_arburst )                             ,
  .m_memory_ar_lock                (mem_core_arlock  )                            ,
  .m_memory_ar_cache               (mem_core_arcache )                             ,
  .m_memory_ar_prot                (mem_core_arprot  )                            ,
  .m_memory_ar_qos                 (mem_core_arqos   )                           ,
  .m_memory_r_ready                (mem_core_rready  )                       ,
  .m_memory_r_valid                (mem_core_rvalid  )                       ,
  .m_memory_r_id                   (mem_core_rid     )                         ,
  .m_memory_r_data                 (mem_core_rdata   )                           ,
  .m_memory_r_resp                 (mem_core_rresp   )                           ,
  .m_memory_r_last                 (mem_core_rlast   )                           ,
  .m_peripheral_aw_ready            (peri_awready  )                            ,
  .m_peripheral_aw_valid            (peri_awvalid  )                            ,
  .m_peripheral_aw_id              (peri_awid     )                              ,
  .m_peripheral_aw_addr            (peri_awaddr   )                                ,
  .m_peripheral_aw_len             (peri_awlen    )                               ,
  .m_peripheral_aw_size            (peri_awsize   )                                ,
  .m_peripheral_aw_burst            (peri_awburst  )                                 ,
  .m_peripheral_aw_lock            (peri_awlock   )                                ,
  .m_peripheral_aw_cache            (peri_awcache  )                                 ,
  .m_peripheral_aw_prot            (peri_awprot   )                                ,
  .m_peripheral_aw_qos             (peri_awqos    )                               ,
  .m_peripheral_w_ready             (peri_wready   )                           ,
  .m_peripheral_w_valid             (peri_wvalid   )                           ,
  .m_peripheral_w_data              (peri_wdata    )                               ,
  .m_peripheral_w_strb              (peri_wstrb    )                               ,
  .m_peripheral_w_last              (peri_wlast    )                               ,
  .m_peripheral_b_ready             (peri_bready   )                           ,
  .m_peripheral_b_valid             (peri_bvalid   )                           ,
  .m_peripheral_b_id                (peri_bid      )                             ,
  .m_peripheral_b_resp              (peri_bresp    )                               ,
  .m_peripheral_ar_ready            (peri_arready  )                            ,
  .m_peripheral_ar_valid            (peri_arvalid  )                            ,
  .m_peripheral_ar_id               (peri_arid     )                              ,
  .m_peripheral_ar_addr             (peri_araddr   )                                ,
  .m_peripheral_ar_len              (peri_arlen    )                               ,
  .m_peripheral_ar_size             (peri_arsize   )                                ,
  .m_peripheral_ar_burst           (peri_arburst  )                                 ,
  .m_peripheral_ar_lock             (peri_arlock   )                                ,
  .m_peripheral_ar_cache            (peri_arcache  )                                 ,
  .m_peripheral_ar_prot             (peri_arprot   )                                ,
  .m_peripheral_ar_qos              (peri_arqos    )                               ,
  .m_peripheral_r_ready             (peri_rready   )                           ,
  .m_peripheral_r_valid             (peri_rvalid   )                           ,
  .m_peripheral_r_id                (peri_rid      )                             ,
  .m_peripheral_r_data              (peri_rdata    )                               ,
  .m_peripheral_r_resp              (peri_rresp    )                               ,
  .m_peripheral_r_last              (peri_rlast    )                               ,
  .s_dma_aw_ready                   (dma_core_awready )                     ,
  .s_dma_aw_valid                   (dma_core_awvalid )                     ,
  .s_dma_aw_id                     (dma_core_awid    )                       ,
  .s_dma_aw_addr                  (dma_core_awaddr[35:0]  )                         ,
  .s_dma_aw_len                    (dma_core_awlen   )                        ,
  .s_dma_aw_size                   (dma_core_awsize  )                         ,
  .s_dma_aw_burst                   (dma_core_awburst )                          ,
  .s_dma_aw_lock                  (dma_core_awlock  )                         ,
  .s_dma_aw_cache                   (dma_core_awcache )                          ,
  .s_dma_aw_prot                   (dma_core_awprot  )                         ,
  .s_dma_aw_qos                    (dma_core_awqos   )                        ,
  .s_dma_w_ready                  (dma_core_wready  )                    ,
  .s_dma_w_valid                   (dma_core_wvalid  )                    ,
  .s_dma_w_data                    (dma_core_wdata   )                        ,
  .s_dma_w_strb                    (dma_core_wstrb   )                        ,
  .s_dma_w_last                   (dma_core_wlast   )                        ,
  .s_dma_b_ready                   (dma_core_bready  )                    ,
  .s_dma_b_valid                  (dma_core_bvalid  )                    ,
  .s_dma_b_id                      (dma_core_bid     )                      ,
  .s_dma_b_resp                    (dma_core_bresp   )                        ,
  .s_dma_ar_ready                   (dma_core_arready )                     ,
  .s_dma_ar_valid                   (dma_core_arvalid )                     ,
  .s_dma_ar_id                     (dma_core_arid    )                       ,
  .s_dma_ar_addr                   (dma_core_araddr[35:0]  )                         ,
  .s_dma_ar_len                    (dma_core_arlen   )                        ,
  .s_dma_ar_size                   (dma_core_arsize  )                         ,
  .s_dma_ar_burst                   (dma_core_arburst )                          ,
  .s_dma_ar_lock                   (dma_core_arlock  )                         ,
  .s_dma_ar_cache                   (dma_core_arcache )                          ,
  .s_dma_ar_prot                   (dma_core_arprot  )                         ,
  .s_dma_ar_qos                    (dma_core_arqos   )                        ,
  .s_dma_r_ready                   (dma_core_rready  )                    ,
  .s_dma_r_valid                   (dma_core_rvalid  )                    ,
  .s_dma_r_id                      (dma_core_rid     )                      ,
  .s_dma_r_data                    (dma_core_rdata   )                        ,
  .s_dma_r_resp                    (dma_core_rresp   )                        ,
  .s_dma_r_last                    (dma_core_rlast   )                        ,
  
  .io_systemjtag_jtag_TCK          (io_systemjtag_jtag_TCK),
  .io_systemjtag_jtag_TMS          (io_systemjtag_jtag_TMS),
  .io_systemjtag_jtag_TDI          (io_systemjtag_jtag_TDI),
  .io_systemjtag_jtag_TDO_data     (io_systemjtag_jtag_TDO_data),
  .io_systemjtag_jtag_TDO_driven   (io_systemjtag_jtag_TDO_driven),
  .io_systemjtag_reset             (io_systemjtag_reset),
  .io_systemjtag_mfr_id            (11'h11),
  .io_systemjtag_part_number       (16'h16),
  .io_systemjtag_version           (4'h4),

  .io_riscv_rst_vec_0              (38'h10000000),
  .dft_lgc_rst_n                   (1'b0),
  .scan_mode                       (1'b0),
  .dft_mode                        (1'b0),
  .rtc_clock                       (rtc_clk),

  .io_clock                        (sys_clk_i/*cpu_clock  */                        ),
  .io_reset                        (~sys_rstn_i/*cpu_global_reset  */                 ),
  .io_extIntrs                     (io_extIntrs  )
);

endmodule
