module XSTop_wrapper(
  input           sys_clk_i,    
  input           sys_rstn_i, 
  input           osc_clock,        //24MHz
  input           outer_clock,      //Max : 2.4GHz
  input           global_reset,     //24MHz

  input  [3:0]    pll_bypass_sel,   //apb clk : 100MHz
  output          pll0_lock,
  output          pll0_clk_div_1024,
  output [11:0]   pll0_test_calout,

  input  [15:0]   soc_to_cpu,   // none
  output [15:0]   cpu_to_soc,   //none

  input  [63:0]   io_extIntrs,   // come from IPs, Max : 600MHz

  input  [15:0]   io_sram_config,  //apb clk : 100MHz

  input           io_systemjtag_jtag_TCK,         // come from gpio
  input           io_systemjtag_jtag_TMS,         // come from gpio
  input           io_systemjtag_jtag_TDI,         // come from gpio
  output          io_systemjtag_jtag_TDO_data,    // come from gpio
  output          io_systemjtag_jtag_TDO_driven,  // come from gpio
  input           io_systemjtag_reset,            // come from gpio

// peri bus   //400MHz
// dma bus    //800MHz
// mem bus    //800MHz

  (*mark_debug="true"*) output          dma_core_awready,
  (*mark_debug="true"*) input           dma_core_awvalid,
  (*mark_debug="true"*) input  [13:0]   dma_core_awid,
  (*mark_debug="true"*) input  [35:0]   dma_core_awaddr,
  (*mark_debug="true"*) input  [7:0]    dma_core_awlen,
  (*mark_debug="true"*) input  [2:0]    dma_core_awsize,
  (*mark_debug="true"*) input  [1:0]    dma_core_awburst,
  (*mark_debug="true"*) input           dma_core_awlock,
  (*mark_debug="true"*) input  [3:0]    dma_core_awcache,
  (*mark_debug="true"*) input  [2:0]    dma_core_awprot,
  (*mark_debug="true"*) input  [3:0]    dma_core_awqos,
  (*mark_debug="true"*) output          dma_core_wready,
  (*mark_debug="true"*) input           dma_core_wvalid,
  (*mark_debug="true"*) input  [255:0]  dma_core_wdata,
  (*mark_debug="true"*) input  [31:0]   dma_core_wstrb,
  (*mark_debug="true"*) input           dma_core_wlast,
  (*mark_debug="true"*) input           dma_core_bready,
  (*mark_debug="true"*) output          dma_core_bvalid,
  (*mark_debug="true"*) output [13:0]   dma_core_bid,
  (*mark_debug="true"*) output [1:0]    dma_core_bresp,
  (*mark_debug="true"*) output          dma_core_arready,
  (*mark_debug="true"*) input           dma_core_arvalid,
  (*mark_debug="true"*) input  [13:0]   dma_core_arid,
  (*mark_debug="true"*) input  [35:0]   dma_core_araddr,
  (*mark_debug="true"*) input  [7:0]    dma_core_arlen,
  (*mark_debug="true"*) input  [2:0]    dma_core_arsize,
  (*mark_debug="true"*) input  [1:0]    dma_core_arburst,
  (*mark_debug="true"*) input           dma_core_arlock,
  (*mark_debug="true"*) input  [3:0]    dma_core_arcache,
  (*mark_debug="true"*) input  [2:0]    dma_core_arprot,
  (*mark_debug="true"*) input  [3:0]    dma_core_arqos,
  (*mark_debug="true"*) input           dma_core_rready,
  (*mark_debug="true"*) output          dma_core_rvalid,
  (*mark_debug="true"*) output [13:0]   dma_core_rid,
  (*mark_debug="true"*) output [255:0]  dma_core_rdata,
  (*mark_debug="true"*) output [1:0]    dma_core_rresp,
  (*mark_debug="true"*) output          dma_core_rlast,
  
  (*mark_debug="true"*) input           peri_awready,
  (*mark_debug="true"*) output          peri_awvalid,
  (*mark_debug="true"*) output [1:0]    peri_awid,
  (*mark_debug="true"*) output [30:0]   peri_awaddr,
  (*mark_debug="true"*) output [7:0]    peri_awlen,
  (*mark_debug="true"*) output [2:0]    peri_awsize,
  (*mark_debug="true"*) output [1:0]    peri_awburst,
  (*mark_debug="true"*) output          peri_awlock,
  (*mark_debug="true"*) output [3:0]    peri_awcache,
  (*mark_debug="true"*) output [2:0]    peri_awprot,
  (*mark_debug="true"*) output [3:0]    peri_awqos,
  (*mark_debug="true"*) input           peri_wready,
  (*mark_debug="true"*) output          peri_wvalid,
  (*mark_debug="true"*) output [63:0]   peri_wdata,
  (*mark_debug="true"*) output [7:0]    peri_wstrb,
  (*mark_debug="true"*) output          peri_wlast,
  (*mark_debug="true"*) output          peri_bready,
  (*mark_debug="true"*) input           peri_bvalid,
  (*mark_debug="true"*) input  [1:0]    peri_bid,
  (*mark_debug="true"*) input  [1:0]    peri_bresp,
  (*mark_debug="true"*) input           peri_arready,
  (*mark_debug="true"*) output          peri_arvalid,
  (*mark_debug="true"*) output [1:0]    peri_arid,
  (*mark_debug="true"*) output [30:0]   peri_araddr,
  (*mark_debug="true"*) output [7:0]    peri_arlen,
  (*mark_debug="true"*) output [2:0]    peri_arsize,
  (*mark_debug="true"*) output [1:0]    peri_arburst,
  (*mark_debug="true"*) output          peri_arlock,
  (*mark_debug="true"*) output [3:0]    peri_arcache,
  (*mark_debug="true"*) output [2:0]    peri_arprot,
  (*mark_debug="true"*) output [3:0]    peri_arqos,
  (*mark_debug="true"*) output          peri_rready,
  (*mark_debug="true"*) input           peri_rvalid,
  (*mark_debug="true"*) input  [1:0]    peri_rid,
  (*mark_debug="true"*) input  [63:0]   peri_rdata,
  (*mark_debug="true"*) input  [1:0]    peri_rresp,
  (*mark_debug="true"*) input           peri_rlast,
  
  (*mark_debug="true"*) input           mem_core_awready,
  (*mark_debug="true"*) output          mem_core_awvalid,
  (*mark_debug="true"*) output [13:0]   mem_core_awid,
  (*mark_debug="true"*) output [35:0]   mem_core_awaddr,
  (*mark_debug="true"*) output [7:0]    mem_core_awlen,
  (*mark_debug="true"*) output [2:0]    mem_core_awsize,
  (*mark_debug="true"*) output [1:0]    mem_core_awburst,
  (*mark_debug="true"*) output          mem_core_awlock,
  (*mark_debug="true"*) output [3:0]    mem_core_awcache,
  (*mark_debug="true"*) output [2:0]    mem_core_awprot,
  (*mark_debug="true"*) output [3:0]    mem_core_awqos,
  (*mark_debug="true"*) input           mem_core_wready,
  (*mark_debug="true"*) output          mem_core_wvalid,
  (*mark_debug="true"*) output [255:0]  mem_core_wdata,
  (*mark_debug="true"*) output [31:0]   mem_core_wstrb,
  (*mark_debug="true"*) output          mem_core_wlast,
  (*mark_debug="true"*) output          mem_core_bready,
  (*mark_debug="true"*) input           mem_core_bvalid,
  (*mark_debug="true"*) input  [13:0]   mem_core_bid,
  (*mark_debug="true"*) input  [1:0]    mem_core_bresp,
  (*mark_debug="true"*) input           mem_core_arready,
  (*mark_debug="true"*) output          mem_core_arvalid,
  (*mark_debug="true"*) output [13:0]   mem_core_arid,
  (*mark_debug="true"*) output [35:0]   mem_core_araddr,
  (*mark_debug="true"*) output [7:0]    mem_core_arlen,
  (*mark_debug="true"*) output [2:0]    mem_core_arsize,
  (*mark_debug="true"*) output [1:0]    mem_core_arburst,
  (*mark_debug="true"*) output          mem_core_arlock,
  (*mark_debug="true"*) output [3:0]    mem_core_arcache,
  (*mark_debug="true"*) output [2:0]    mem_core_arprot,
  (*mark_debug="true"*) output [3:0]    mem_core_arqos,
  (*mark_debug="true"*) output          mem_core_rready,
  (*mark_debug="true"*) input           mem_core_rvalid,
  (*mark_debug="true"*) input  [13:0]   mem_core_rid,
  (*mark_debug="true"*) input  [255:0]  mem_core_rdata,
  (*mark_debug="true"*) input  [1:0]    mem_core_rresp,
  (*mark_debug="true"*) input           mem_core_rlast
);

  wire          cpu_clock       ;
  wire          cpu_global_reset;
  wire          global_reset_sync;

  wire [31:0]   pll0_config_0;
  wire [31:0]   pll0_config_1;
  wire [31:0]   pll0_config_2;
  wire [31:0]   pll0_config_3;
  wire [31:0]   pll0_config_4;
  wire [31:0]   pll0_config_5;
//  wire [31:0]   pll0_config_5 = 32'h3;

assign cpu_to_soc = 32'h0;


XSTop  u_XSTop(
  .memory_0_awready                (mem_core_awready )                        ,
  .memory_0_awvalid                (mem_core_awvalid )                        ,
  .memory_0_awid                   (mem_core_awid    )                          ,
  .memory_0_awaddr                 (mem_core_awaddr  )                            ,
  .memory_0_awlen                  (mem_core_awlen   )                           ,
  .memory_0_awsize                 (mem_core_awsize  )                            ,
  .memory_0_awburst                (mem_core_awburst )                             ,
  .memory_0_awlock                 (mem_core_awlock  )                            ,
  .memory_0_awcache                (mem_core_awcache )                             ,
  .memory_0_awprot                 (mem_core_awprot  )                            ,
  .memory_0_awqos                  (mem_core_awqos   )                           ,
  .memory_0_wready                 (mem_core_wready  )                       ,
  .memory_0_wvalid                 (mem_core_wvalid  )                       ,
  .memory_0_wdata                  (mem_core_wdata   )                           ,
  .memory_0_wstrb                  (mem_core_wstrb   )                           ,
  .memory_0_wlast                  (mem_core_wlast   )                           ,
  .memory_0_bready                 (mem_core_bready  )                       ,
  .memory_0_bvalid                 (mem_core_bvalid  )                       ,
  .memory_0_bid                    (mem_core_bid     )                         ,
  .memory_0_bresp                  (mem_core_bresp   )                           ,
  .memory_0_arready                (mem_core_arready )                        ,
  .memory_0_arvalid                (mem_core_arvalid )                        ,
  .memory_0_arid                   (mem_core_arid    )                          ,
  .memory_0_araddr                 (mem_core_araddr  )                            ,
  .memory_0_arlen                  (mem_core_arlen   )                           ,
  .memory_0_arsize                 (mem_core_arsize  )                            ,
  .memory_0_arburst                (mem_core_arburst )                             ,
  .memory_0_arlock                 (mem_core_arlock  )                            ,
  .memory_0_arcache                (mem_core_arcache )                             ,
  .memory_0_arprot                 (mem_core_arprot  )                            ,
  .memory_0_arqos                  (mem_core_arqos   )                           ,
  .memory_0_rready                 (mem_core_rready  )                       ,
  .memory_0_rvalid                 (mem_core_rvalid  )                       ,
  .memory_0_rid                    (mem_core_rid     )                         ,
  .memory_0_rdata                  (mem_core_rdata   )                           ,
  .memory_0_rresp                  (mem_core_rresp   )                           ,
  .memory_0_rlast                  (mem_core_rlast   )                           ,
  .peripheral_0_awready            (peri_awready  )                            ,
  .peripheral_0_awvalid            (peri_awvalid  )                            ,
  .peripheral_0_awid               (peri_awid     )                              ,
  .peripheral_0_awaddr             (peri_awaddr   )                                ,
  .peripheral_0_awlen              (peri_awlen    )                               ,
  .peripheral_0_awsize             (peri_awsize   )                                ,
  .peripheral_0_awburst            (peri_awburst  )                                 ,
  .peripheral_0_awlock             (peri_awlock   )                                ,
  .peripheral_0_awcache            (peri_awcache  )                                 ,
  .peripheral_0_awprot             (peri_awprot   )                                ,
  .peripheral_0_awqos              (peri_awqos    )                               ,
  .peripheral_0_wready             (peri_wready   )                           ,
  .peripheral_0_wvalid             (peri_wvalid   )                           ,
  .peripheral_0_wdata              (peri_wdata    )                               ,
  .peripheral_0_wstrb              (peri_wstrb    )                               ,
  .peripheral_0_wlast              (peri_wlast    )                               ,
  .peripheral_0_bready             (peri_bready   )                           ,
  .peripheral_0_bvalid             (peri_bvalid   )                           ,
  .peripheral_0_bid                (peri_bid      )                             ,
  .peripheral_0_bresp              (peri_bresp    )                               ,
  .peripheral_0_arready            (peri_arready  )                            ,
  .peripheral_0_arvalid            (peri_arvalid  )                            ,
  .peripheral_0_arid               (peri_arid     )                              ,
  .peripheral_0_araddr             (peri_araddr   )                                ,
  .peripheral_0_arlen              (peri_arlen    )                               ,
  .peripheral_0_arsize             (peri_arsize   )                                ,
  .peripheral_0_arburst            (peri_arburst  )                                 ,
  .peripheral_0_arlock             (peri_arlock   )                                ,
  .peripheral_0_arcache            (peri_arcache  )                                 ,
  .peripheral_0_arprot             (peri_arprot   )                                ,
  .peripheral_0_arqos              (peri_arqos    )                               ,
  .peripheral_0_rready             (peri_rready   )                           ,
  .peripheral_0_rvalid             (peri_rvalid   )                           ,
  .peripheral_0_rid                (peri_rid      )                             ,
  .peripheral_0_rdata              (peri_rdata    )                               ,
  .peripheral_0_rresp              (peri_rresp    )                               ,
  .peripheral_0_rlast              (peri_rlast    )                               ,
  .dma_0_awready                   (dma_core_awready )                     ,
  .dma_0_awvalid                   (dma_core_awvalid )                     ,
  .dma_0_awid                      (dma_core_awid    )                       ,
  .dma_0_awaddr                    (dma_core_awaddr[35:0]  )                         ,
  .dma_0_awlen                     (dma_core_awlen   )                        ,
  .dma_0_awsize                    (dma_core_awsize  )                         ,
  .dma_0_awburst                   (dma_core_awburst )                          ,
  .dma_0_awlock                    (dma_core_awlock  )                         ,
  .dma_0_awcache                   (dma_core_awcache )                          ,
  .dma_0_awprot                    (dma_core_awprot  )                         ,
  .dma_0_awqos                     (dma_core_awqos   )                        ,
  .dma_0_wready                    (dma_core_wready  )                    ,
  .dma_0_wvalid                    (dma_core_wvalid  )                    ,
  .dma_0_wdata                     (dma_core_wdata   )                        ,
  .dma_0_wstrb                     (dma_core_wstrb   )                        ,
  .dma_0_wlast                     (dma_core_wlast   )                        ,
  .dma_0_bready                    (dma_core_bready  )                    ,
  .dma_0_bvalid                    (dma_core_bvalid  )                    ,
  .dma_0_bid                       (dma_core_bid     )                      ,
  .dma_0_bresp                     (dma_core_bresp   )                        ,
  .dma_0_arready                   (dma_core_arready )                     ,
  .dma_0_arvalid                   (dma_core_arvalid )                     ,
  .dma_0_arid                      (dma_core_arid    )                       ,
  .dma_0_araddr                    (dma_core_araddr[35:0]  )                         ,
  .dma_0_arlen                     (dma_core_arlen   )                        ,
  .dma_0_arsize                    (dma_core_arsize  )                         ,
  .dma_0_arburst                   (dma_core_arburst )                          ,
  .dma_0_arlock                    (dma_core_arlock  )                         ,
  .dma_0_arcache                   (dma_core_arcache )                          ,
  .dma_0_arprot                    (dma_core_arprot  )                         ,
  .dma_0_arqos                     (dma_core_arqos   )                        ,
  .dma_0_rready                    (dma_core_rready  )                    ,
  .dma_0_rvalid                    (dma_core_rvalid  )                    ,
  .dma_0_rid                       (dma_core_rid     )                      ,
  .dma_0_rdata                     (dma_core_rdata   )                        ,
  .dma_0_rresp                     (dma_core_rresp   )                        ,
  .dma_0_rlast                     (dma_core_rlast   )                        ,
  
  .io_systemjtag_jtag_TCK          (io_systemjtag_jtag_TCK),
  .io_systemjtag_jtag_TMS          (io_systemjtag_jtag_TMS),
  .io_systemjtag_jtag_TDI          (io_systemjtag_jtag_TDI),
  .io_systemjtag_jtag_TDO_data     (io_systemjtag_jtag_TDO_data),
  .io_systemjtag_jtag_TDO_driven   (io_systemjtag_jtag_TDO_driven),
  .io_systemjtag_reset             (io_systemjtag_reset),
  .io_systemjtag_mfr_id            (11'h11),
  .io_systemjtag_part_number       (16'h16),
  .io_systemjtag_version           (4'h4),

  .io_clock                        (sys_clk_i/*cpu_clock  */                        ),
  .io_reset                        (~sys_rstn_i/*cpu_global_reset  */                 ),
  .io_extIntrs                     (io_extIntrs  )
);

endmodule
