`include "DSEMacro.v"

module XSTop_wrapper_dse(
  input           clock,
  input           reset,

  output [63:0]   io_extIntrs,
  output          out_enable,
  output [`DEG_DATA_WIDTH+`MAGIC_NUM_WIDTH-1:0] out_io_data,

  output          dma_core_awready,
  input           dma_core_awvalid,
  input  [13:0]   dma_core_awid,
  input  [35:0]   dma_core_awaddr,
  input  [7:0]    dma_core_awlen,
  input  [2:0]    dma_core_awsize,
  input  [1:0]    dma_core_awburst,
  input           dma_core_awlock,
  input  [3:0]    dma_core_awcache,
  input  [2:0]    dma_core_awprot,
  input  [3:0]    dma_core_awqos,
  output          dma_core_wready,
  input           dma_core_wvalid,
  input  [255:0]  dma_core_wdata,
  input  [31:0]   dma_core_wstrb,
  input           dma_core_wlast,
  input           dma_core_bready,
  output          dma_core_bvalid,
  output [13:0]   dma_core_bid,
  output [1:0]    dma_core_bresp,
  output          dma_core_arready,
  input           dma_core_arvalid,
  input  [13:0]   dma_core_arid,
  input  [35:0]   dma_core_araddr,
  input  [7:0]    dma_core_arlen,
  input  [2:0]    dma_core_arsize,
  input  [1:0]    dma_core_arburst,
  input           dma_core_arlock,
  input  [3:0]    dma_core_arcache,
  input  [2:0]    dma_core_arprot,
  input  [3:0]    dma_core_arqos,
  input           dma_core_rready,
  output          dma_core_rvalid,
  output [13:0]   dma_core_rid,
  output [255:0]  dma_core_rdata,
  output [1:0]    dma_core_rresp,
  output          dma_core_rlast,
  
  input           peri_awready,
  output          peri_awvalid,
  output [1:0]    peri_awid,
  output [30:0]   peri_awaddr,
  output [7:0]    peri_awlen,
  output [2:0]    peri_awsize,
  output [1:0]    peri_awburst,
  output          peri_awlock,
  output [3:0]    peri_awcache,
  output [2:0]    peri_awprot,
  output [3:0]    peri_awqos,
  input           peri_wready,
  output          peri_wvalid,
  output [63:0]   peri_wdata,
  output [7:0]    peri_wstrb,
  output          peri_wlast,
  output          peri_bready,
  input           peri_bvalid,
  input  [1:0]    peri_bid,
  input  [1:0]    peri_bresp,
  input           peri_arready,
  output          peri_arvalid,
  output [1:0]    peri_arid,
  output [30:0]   peri_araddr,
  output [7:0]    peri_arlen,
  output [2:0]    peri_arsize,
  output [1:0]    peri_arburst,
  output          peri_arlock,
  output [3:0]    peri_arcache,
  output [2:0]    peri_arprot,
  output [3:0]    peri_arqos,
  output          peri_rready,
  input           peri_rvalid,
  input  [1:0]    peri_rid,
  input  [63:0]   peri_rdata,
  input  [1:0]    peri_rresp,
  input           peri_rlast,
  
  input           mem_core_awready,
  output          mem_core_awvalid,
  output [13:0]   mem_core_awid,
  output [35:0]   mem_core_awaddr,
  output [7:0]    mem_core_awlen,
  output [2:0]    mem_core_awsize,
  output [1:0]    mem_core_awburst,
  output          mem_core_awlock,
  output [3:0]    mem_core_awcache,
  output [2:0]    mem_core_awprot,
  output [3:0]    mem_core_awqos,
  input           mem_core_wready,
  output          mem_core_wvalid,
  output [255:0]  mem_core_wdata,
  output [31:0]   mem_core_wstrb,
  output          mem_core_wlast,
  output          mem_core_bready,
  input           mem_core_bvalid,
  input  [13:0]   mem_core_bid,
  input  [1:0]    mem_core_bresp,
  input           mem_core_arready,
  output          mem_core_arvalid,
  output [13:0]   mem_core_arid,
  output [35:0]   mem_core_araddr,
  output [7:0]    mem_core_arlen,
  output [2:0]    mem_core_arsize,
  output [1:0]    mem_core_arburst,
  output          mem_core_arlock,
  output [3:0]    mem_core_arcache,
  output [2:0]    mem_core_arprot,
  output [3:0]    mem_core_arqos,
  output          mem_core_rready,
  input           mem_core_rvalid,
  input  [13:0]   mem_core_rid,
  input  [255:0]  mem_core_rdata,
  input  [1:0]    mem_core_rresp,
  input           mem_core_rlast
);

  wire dse_reset_valid;
  wire [35:0] dse_reset_vector;
  wire [63:0] dse_epoch;

  // define performance counter wires
  wire deg_out_enable;
  wire [5:0] deg_valids;
  wire [`DEG_DATA_WIDTH-1:0] deg_out_data;  // [16000:0] is valid data
  wire [`PERF_DATA_WIDTH-1:0] perf_out_data;
  wire dse_endpoint_out_enable;
  wire [`DEG_DATA_WIDTH+`MAGIC_NUM_WIDTH-1:0] dse_endpoint_out_data;

  XSTop  u_XSTop(
    .memory_0_awready                (mem_core_awready )                        ,
    .memory_0_awvalid                (mem_core_awvalid )                        ,
    .memory_0_awid                   (mem_core_awid    )                          ,
    .memory_0_awaddr                 (mem_core_awaddr  )                            ,
    .memory_0_awlen                  (mem_core_awlen   )                           ,
    .memory_0_awsize                 (mem_core_awsize  )                            ,
    .memory_0_awburst                (mem_core_awburst )                             ,
    .memory_0_awlock                 (mem_core_awlock  )                            ,
    .memory_0_awcache                (mem_core_awcache )                             ,
    .memory_0_awprot                 (mem_core_awprot  )                            ,
    .memory_0_awqos                  (mem_core_awqos   )                           ,
    .memory_0_wready                 (mem_core_wready  )                       ,
    .memory_0_wvalid                 (mem_core_wvalid  )                       ,
    .memory_0_wdata                  (mem_core_wdata   )                           ,
    .memory_0_wstrb                  (mem_core_wstrb   )                           ,
    .memory_0_wlast                  (mem_core_wlast   )                           ,
    .memory_0_bready                 (mem_core_bready  )                       ,
    .memory_0_bvalid                 (mem_core_bvalid  )                       ,
    .memory_0_bid                    (mem_core_bid     )                         ,
    .memory_0_bresp                  (mem_core_bresp   )                           ,
    .memory_0_arready                (mem_core_arready )                        ,
    .memory_0_arvalid                (mem_core_arvalid )                        ,
    .memory_0_arid                   (mem_core_arid    )                          ,
    .memory_0_araddr                 (mem_core_araddr  )                            ,
    .memory_0_arlen                  (mem_core_arlen   )                           ,
    .memory_0_arsize                 (mem_core_arsize  )                            ,
    .memory_0_arburst                (mem_core_arburst )                             ,
    .memory_0_arlock                 (mem_core_arlock  )                            ,
    .memory_0_arcache                (mem_core_arcache )                             ,
    .memory_0_arprot                 (mem_core_arprot  )                            ,
    .memory_0_arqos                  (mem_core_arqos   )                           ,
    .memory_0_rready                 (mem_core_rready  )                       ,
    .memory_0_rvalid                 (mem_core_rvalid  )                       ,
    .memory_0_rid                    (mem_core_rid     )                         ,
    .memory_0_rdata                  (mem_core_rdata   )                           ,
    .memory_0_rresp                  (mem_core_rresp   )                           ,
    .memory_0_rlast                  (mem_core_rlast   )                           ,
    .peripheral_0_awready            (peri_awready  )                            ,
    .peripheral_0_awvalid            (peri_awvalid  )                            ,
    .peripheral_0_awid               (peri_awid     )                              ,
    .peripheral_0_awaddr             (peri_awaddr   )                                ,
    .peripheral_0_awlen              (peri_awlen    )                               ,
    .peripheral_0_awsize             (peri_awsize   )                                ,
    .peripheral_0_awburst            (peri_awburst  )                                 ,
    .peripheral_0_awlock             (peri_awlock   )                                ,
    .peripheral_0_awcache            (peri_awcache  )                                 ,
    .peripheral_0_awprot             (peri_awprot   )                                ,
    .peripheral_0_awqos              (peri_awqos    )                               ,
    .peripheral_0_wready             (peri_wready   )                           ,
    .peripheral_0_wvalid             (peri_wvalid   )                           ,
    .peripheral_0_wdata              (peri_wdata    )                               ,
    .peripheral_0_wstrb              (peri_wstrb    )                               ,
    .peripheral_0_wlast              (peri_wlast    )                               ,
    .peripheral_0_bready             (peri_bready   )                           ,
    .peripheral_0_bvalid             (peri_bvalid   )                           ,
    .peripheral_0_bid                (peri_bid      )                             ,
    .peripheral_0_bresp              (peri_bresp    )                               ,
    .peripheral_0_arready            (peri_arready  )                            ,
    .peripheral_0_arvalid            (peri_arvalid  )                            ,
    .peripheral_0_arid               (peri_arid     )                              ,
    .peripheral_0_araddr             (peri_araddr   )                                ,
    .peripheral_0_arlen              (peri_arlen    )                               ,
    .peripheral_0_arsize             (peri_arsize   )                                ,
    .peripheral_0_arburst            (peri_arburst  )                                 ,
    .peripheral_0_arlock             (peri_arlock   )                                ,
    .peripheral_0_arcache            (peri_arcache  )                                 ,
    .peripheral_0_arprot             (peri_arprot   )                                ,
    .peripheral_0_arqos              (peri_arqos    )                               ,
    .peripheral_0_rready             (peri_rready   )                           ,
    .peripheral_0_rvalid             (peri_rvalid   )                           ,
    .peripheral_0_rid                (peri_rid      )                             ,
    .peripheral_0_rdata              (peri_rdata    )                               ,
    .peripheral_0_rresp              (peri_rresp    )                               ,
    .peripheral_0_rlast              (peri_rlast    )                               ,
    .dma_0_awready                   (dma_core_awready )                     ,
    .dma_0_awvalid                   (dma_core_awvalid )                     ,
    .dma_0_awid                      (dma_core_awid    )                       ,
    .dma_0_awaddr                    (dma_core_awaddr[35:0]  )                         ,
    .dma_0_awlen                     (dma_core_awlen   )                        ,
    .dma_0_awsize                    (dma_core_awsize  )                         ,
    .dma_0_awburst                   (dma_core_awburst )                          ,
    .dma_0_awlock                    (dma_core_awlock  )                         ,
    .dma_0_awcache                   (dma_core_awcache )                          ,
    .dma_0_awprot                    (dma_core_awprot  )                         ,
    .dma_0_awqos                     (dma_core_awqos   )                        ,
    .dma_0_wready                    (dma_core_wready  )                    ,
    .dma_0_wvalid                    (dma_core_wvalid  )                    ,
    .dma_0_wdata                     (dma_core_wdata   )                        ,
    .dma_0_wstrb                     (dma_core_wstrb   )                        ,
    .dma_0_wlast                     (dma_core_wlast   )                        ,
    .dma_0_bready                    (dma_core_bready  )                    ,
    .dma_0_bvalid                    (dma_core_bvalid  )                    ,
    .dma_0_bid                       (dma_core_bid     )                      ,
    .dma_0_bresp                     (dma_core_bresp   )                        ,
    .dma_0_arready                   (dma_core_arready )                     ,
    .dma_0_arvalid                   (dma_core_arvalid )                     ,
    .dma_0_arid                      (dma_core_arid    )                       ,
    .dma_0_araddr                    (dma_core_araddr[35:0]  )                         ,
    .dma_0_arlen                     (dma_core_arlen   )                        ,
    .dma_0_arsize                    (dma_core_arsize  )                         ,
    .dma_0_arburst                   (dma_core_arburst )                          ,
    .dma_0_arlock                    (dma_core_arlock  )                         ,
    .dma_0_arcache                   (dma_core_arcache )                          ,
    .dma_0_arprot                    (dma_core_arprot  )                         ,
    .dma_0_arqos                     (dma_core_arqos   )                        ,
    .dma_0_rready                    (dma_core_rready  )                    ,
    .dma_0_rvalid                    (dma_core_rvalid  )                    ,
    .dma_0_rid                       (dma_core_rid     )                      ,
    .dma_0_rdata                     (dma_core_rdata   )                        ,
    .dma_0_rresp                     (dma_core_rresp   )                        ,
    .dma_0_rlast                     (dma_core_rlast   )                        ,
    
    .io_systemjtag_jtag_TCK          (_jtag_jtag_TCK),
    .io_systemjtag_jtag_TMS          (_jtag_jtag_TMS),
    .io_systemjtag_jtag_TDI          (_jtag_jtag_TDI),
    .io_systemjtag_jtag_TDO_data     (_l_soc_io_systemjtag_jtag_TDO_data),
    .io_systemjtag_jtag_TDO_driven   (_l_soc_io_systemjtag_jtag_TDO_driven),
    .io_systemjtag_reset             (reset),
    .io_systemjtag_mfr_id            (11'h11),
    .io_systemjtag_part_number       (16'h16),
    .io_systemjtag_version           (4'h4),

    .io_clock                        (clock    ),
    .io_reset                        (reset  ),
    .io_extIntrs                     (io_extIntrs  ),

    .io_instrCnt                        (/* unused */),
    .io_dse_rst                         (reset),
    .io_reset_vector                    (36'h10000000),
    .io_dse_reset_valid                 (dse_reset_valid),
    .io_dse_reset_vec                   (dse_reset_vector),
    .io_dse_max_epoch                   (/* unused */),
    .io_dse_epoch                       (dse_epoch),
    .io_dse_max_instr                   (),
    .deg_out_enable                     (deg_out_enable),
    .deg_out_data                       (deg_out_data),
    .perf_out_data                      (perf_out_data),
    .deg_valids                         (deg_valids)
  );

  SimJTAG #(
    .TICK_DELAY(3)
  ) jtag (	// src/test/scala/top/SimTop.scala:63:20
    .clock           (clock),
    .reset           (reset),
    .jtag_TRSTn      (/* unused */),
    .jtag_TCK        (_jtag_jtag_TCK),
    .jtag_TMS        (_jtag_jtag_TMS),
    .jtag_TDI        (_jtag_jtag_TDI),
    .jtag_TDO_data   (_l_soc_io_systemjtag_jtag_TDO_data),	// src/test/scala/top/SimTop.scala:36:19
    .jtag_TDO_driven (_l_soc_io_systemjtag_jtag_TDO_driven),	// src/test/scala/top/SimTop.scala:36:19
    .enable          (1'h1),	// src/test/scala/top/SimTop.scala:59:20
    .init_done       (~reset),	// src/test/scala/top/SimTop.scala:64:61
    .exit            (/* unused */)
  );

  DSEEndpoint dseendpoint (
    .clock              (clock           ),
    .reset              (reset           ),
    .dse_reset_valid    (dse_reset_valid ),
    .dse_reset_vector   (dse_reset_vector),
    .dse_epoch          (dse_epoch       ),
    .deg_out_enable     (deg_out_enable  ),
    .deg_valids         (deg_valids      ),
    .deg_out_data       (deg_out_data    ),
    .perf_out_data      (perf_out_data   ),
    .out_enable         (dse_endpoint_out_enable),
    .out_data           (dse_endpoint_out_data)
  );

  assign out_enable = dse_endpoint_out_enable;
  assign out_io_data = dse_endpoint_out_data;

endmodule
